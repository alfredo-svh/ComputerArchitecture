module im(clk, addr, IOut);
    //create the array of instructions (size 256, each of 32 bits)
    wire [31:0] inst[260:0];
    
    //initialize variables
    input clk;
    input [31:0] addr;
    output reg [31:0] IOut;
    
    // instructions for the MAX function
        assign inst[0] = 32'b11100010100010110000000000000000;
        assign inst[1] = 32'b11110100100000000101100000000000;
        assign inst[2] = 32'b11110011010000000000000000000000;
        assign inst[3] = 32'b01010011100011100000000000000000;
        assign inst[4] = 32'b00000000000000000000000000000000;
        assign inst[5] = 32'b00000000000000000000000000000000;
        assign inst[6] = 32'b01110011110011000011100000000000;
        assign inst[7] = 32'b10010000000100100000000000000000;
        assign inst[8] = 32'b00000000000000000000000000000000;
        assign inst[9] = 32'b00000000000000000000000000000000;
        assign inst[10] = 32'b01000011110010110011100000000000;
        assign inst[11] = 32'b00000000000000000000000000000000;
        assign inst[12] = 32'b00000000000000000000000000000000;
        assign inst[13] = 32'b11100100010011110000000000000000;
        assign inst[14] = 32'b00000000000000000000000000000000;
        assign inst[15] = 32'b00000000000000000000000000000000;
        assign inst[16] = 32'b01110101000100010010100000000000;
        assign inst[17] = 32'b10110000000011010000000000000000;
        assign inst[18] = 32'b00000000000000000000000000000000;
        assign inst[19] = 32'b00000000000000000000000000000000;
        assign inst[20] = 32'b00000000000000000000000000000000;
        assign inst[21] = 32'b01000010100000000100010000000000;
        assign inst[22] = 32'b10000000000011010000000000000000;
        assign inst[23] = 32'b00000000000000000000000000000000;
        assign inst[24] = 32'b00000000000000000000000000000000;
    
    
    // instructions for the demo
//    assign inst[0] = 32'b11110000010001000000000000000000;
//    assign inst[1] = 32'b01010000100000010000000000000000;
//    assign inst[2] = 32'b01100000110000010000000000000000;
//    assign inst[3] = 32'b11110010100000000010010000000000;
//    assign inst[4] = 32'b00000000000000000000000000000000;
//    assign inst[5] = 32'b00000000000000000000000000000000;
//    assign inst[6] = 32'b10110000000010100000000000000000;
//    assign inst[7] = 32'b00000000000000000000000000000000;
//    assign inst[8] = 32'b00000000000000000000000000000000;
//    assign inst[9] = 32'b00000000000000000000000000000000;
//    assign inst[10] = 32'b00000000000000000000000000000000;
//    assign inst[11] = 32'b01010000100000100000000000000000;
//    assign inst[12] = 32'b00110000000000010000010000000000;
//    assign inst[13] = 32'b11100001000000010000000000000000;
//    assign inst[14] = 32'b01000001010000010000100000000000;
//    assign inst[15] = 32'b00000000000000000000000000000000;
//    assign inst[16] = 32'b01110001100001000000010000000000;
//    assign inst[17] = 32'b11110010110000000010010000000000;
//    assign inst[18] = 32'b00000000000000000000000000000000;
//    assign inst[19] = 32'b00000000000000000000000000000000;
//    assign inst[20] = 32'b10010000000010110000000000000000;
//    assign inst[21] = 32'b00000000000000000000000000000000;
//    assign inst[22] = 32'b00000000000000000000000000000000;
//    assign inst[23] = 32'b00000000000000000000000000000000;
//    assign inst[24] = 32'b00000000000000000000000000000000;
//    assign inst[25] = 32'b01010000100000100000000000000000;
//    assign inst[26] = 32'b10100000000000010000000000000000;
//    assign inst[27] = 32'b00000000000000000000000000000000;
//    assign inst[28] = 32'b00000000000000000000000000000000;
//    assign inst[29] = 32'b00000000000000000000000000000000;
//    assign inst[30] = 32'b00000000000000000000000000000000;    
    
//    assign inst[256] = 32'b10000000000000010000000000000000;
//    assign inst[257] = 32'b00000000000000000000000000000000;
//    assign inst[258] = 32'b00000000000000000000000000000000;
//    assign inst[259] = 32'b00000000000000000000000000000000;
    
    //output the instruction saved at the address taken as input at every positive edge of clock
    always@(negedge clk)
    begin
        IOut = inst[addr];
    end

endmodule